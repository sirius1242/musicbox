`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/23 11:16:25
// Design Name: 
// Module Name: regfile
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module regfile(
    input clk, 
		input rst_n, 
		input [15:0] addr_a, 
		input [15:0] addr_b, 
		input [15:0] addr_c, 
		input [11:0] data_c, 
		input wen_c,
		output wire [11:0] q_a, 
		output wire [11:0] q_b
	);
	integer i;
	reg [11:0] data [0:256];
	always@(posedge clk or negedge rst_n)
	begin
		if (~rst_n)
		begin
			data[0][11:8]<=0;data[0][7:5]<=2;data[0][4:0]<=4;
			data[1][11:8]<=0;data[1][7:5]<=2;data[1][4:0]<=4;
			data[2][11:8]<=0;data[2][7:5]<=2;data[2][4:0]<=4;
			data[3][11:8]<=6;data[3][7:5]<=2;data[3][4:0]<=4;
			data[4][11:8]<=9;data[4][7:5]<=2;data[4][4:0]<=6;
			data[5][11:8]<=9;data[5][7:5]<=2;data[5][4:0]<=2;
			data[6][11:8]<=7;data[6][7:5]<=2;data[6][4:0]<=4;
			data[7][11:8]<=6;data[7][7:5]<=2;data[7][4:0]<=4;
			data[8][11:8]<=4;data[8][7:5]<=2;data[8][4:0]<=6;
			data[9][11:8]<=6;data[9][7:5]<=2;data[9][4:0]<=2;
			data[10][11:8]<=7;data[10][7:5]<=2;data[10][4:0]<=6;
			data[11][11:8]<=7;data[11][7:5]<=2;data[11][4:0]<=2;
			data[12][11:8]<=6;data[12][7:5]<=2;data[12][4:0]<=6;
			data[13][11:8]<=6;data[13][7:5]<=2;data[13][4:0]<=2;
			data[14][11:8]<=4;data[14][7:5]<=2;data[14][4:0]<=6;
			data[15][11:8]<=4;data[15][7:5]<=2;data[15][4:0]<=2;
			data[16][11:8]<=2;data[16][7:5]<=2;data[16][4:0]<=12;
			data[17][11:8]<=9;data[17][7:5]<=2;data[17][4:0]<=4;
			data[18][11:8]<=2;data[18][7:5]<=1;data[18][4:0]<=6;
			data[19][11:8]<=13;data[19][7:5]<=2;data[19][4:0]<=2;
			data[20][11:8]<=4;data[20][7:5]<=1;data[20][4:0]<=2;
			data[21][11:8]<=2;data[21][7:5]<=1;data[21][4:0]<=2;
			data[22][11:8]<=9;data[22][7:5]<=2;data[22][4:0]<=2;
			data[23][11:8]<=6;data[23][7:5]<=2;data[23][4:0]<=2;
			data[24][11:8]<=11;data[24][7:5]<=2;data[24][4:0]<=8;
			data[25][11:8]<=7;data[25][7:5]<=2;data[25][4:0]<=4;
			data[26][11:8]<=0;data[26][7:5]<=2;data[26][4:0]<=2;
			data[27][11:8]<=11;data[27][7:5]<=2;data[27][4:0]<=2;
			data[28][11:8]<=4;data[28][7:5]<=1;data[28][4:0]<=6;
			data[29][11:8]<=2;data[29][7:5]<=2;data[29][4:0]<=4;
			data[30][11:8]<=13;data[30][7:5]<=2;data[30][4:0]<=2;
			data[31][11:8]<=11;data[31][7:5]<=2;data[31][4:0]<=2;
			data[32][11:8]<=9;data[32][7:5]<=2;data[32][4:0]<=2;
			data[33][11:8]<=7;data[33][7:5]<=2;data[33][4:0]<=2;
			data[34][11:8]<=6;data[34][7:5]<=2;data[34][4:0]<=12;
			data[35][11:8]<=9;data[35][7:5]<=2;data[35][4:0]<=2;
			data[36][11:8]<=2;data[36][7:5]<=1;data[36][4:0]<=6;
			data[37][11:8]<=13;data[37][7:5]<=2;data[37][4:0]<=2;
			data[38][11:8]<=4;data[38][7:5]<=1;data[38][4:0]<=2;
			data[39][11:8]<=2;data[39][7:5]<=1;data[39][4:0]<=2;
			data[40][11:8]<=9;data[40][7:5]<=2;data[40][4:0]<=2;
			data[41][11:8]<=6;data[41][7:5]<=2;data[41][4:0]<=2;
			data[42][11:8]<=11;data[42][7:5]<=2;data[42][4:0]<=8;
			data[43][11:8]<=7;data[43][7:5]<=2;data[43][4:0]<=2;
			data[44][11:8]<=11;data[44][7:5]<=2;data[44][4:0]<=2;
			data[45][11:8]<=4;data[45][7:5]<=1;data[45][4:0]<=2;
			data[46][11:8]<=2;data[46][7:5]<=1;data[46][4:0]<=2;
			data[47][11:8]<=13;data[47][7:5]<=2;data[47][4:0]<=4;
			data[48][11:8]<=4;data[48][7:5]<=1;data[48][4:0]<=4;
			data[49][11:8]<=7;data[49][7:5]<=1;data[49][4:0]<=4;
			data[50][11:8]<=13;data[50][7:5]<=2;data[50][4:0]<=4;
			data[51][11:8]<=2;data[51][7:5]<=1;data[51][4:0]<=8;
			data[52][11:8]<=2;data[52][7:5]<=1;data[52][4:0]<=2;
			data[53][11:8]<=0;data[53][7:5]<=2;data[53][4:0]<=2;
			data[54][11:8]<=6;data[54][7:5]<=1;data[54][4:0]<=2;
			data[55][11:8]<=4;data[55][7:5]<=1;data[55][4:0]<=2;
			data[56][11:8]<=13;data[56][7:5]<=2;data[56][4:0]<=8;
			data[57][11:8]<=11;data[57][7:5]<=2;data[57][4:0]<=2;
			data[58][11:8]<=13;data[58][7:5]<=2;data[58][4:0]<=2;
			data[59][11:8]<=2;data[59][7:5]<=1;data[59][4:0]<=2;
			data[60][11:8]<=11;data[60][7:5]<=2;data[60][4:0]<=2;
			data[61][11:8]<=13;data[61][7:5]<=2;data[61][4:0]<=8;
			data[62][11:8]<=9;data[62][7:5]<=2;data[62][4:0]<=2;
			data[63][11:8]<=9;data[63][7:5]<=2;data[63][4:0]<=2;
			data[64][11:8]<=8;data[64][7:5]<=2;data[64][4:0]<=2;
			data[65][11:8]<=9;data[65][7:5]<=2;data[65][4:0]<=2;
			data[66][11:8]<=11;data[66][7:5]<=2;data[66][4:0]<=6;
			data[67][11:8]<=11;data[67][7:5]<=2;data[67][4:0]<=2;
			data[68][11:8]<=4;data[68][7:5]<=1;data[68][4:0]<=4;
			data[69][11:8]<=2;data[69][7:5]<=1;data[69][4:0]<=2;
			data[70][11:8]<=13;data[70][7:5]<=2;data[70][4:0]<=8;
			data[71][11:8]<=13;data[71][7:5]<=2;data[71][4:0]<=2;
			data[72][11:8]<=0;data[72][7:5]<=2;data[72][4:0]<=2;
			data[73][11:8]<=4;data[73][7:5]<=1;data[73][4:0]<=4;
			data[74][11:8]<=4;data[74][7:5]<=1;data[74][4:0]<=6;
			data[75][11:8]<=13;data[75][7:5]<=2;data[75][4:0]<=2;
			data[76][11:8]<=9;data[76][7:5]<=2;data[76][4:0]<=2;
			data[77][11:8]<=9;data[77][7:5]<=2;data[77][4:0]<=2;
			data[78][11:8]<=8;data[78][7:5]<=2;data[78][4:0]<=2;
			data[79][11:8]<=9;data[79][7:5]<=2;data[79][4:0]<=2;
			data[80][11:8]<=6;data[80][7:5]<=1;data[80][4:0]<=8;
			data[81][11:8]<=2;data[81][7:5]<=1;data[81][4:0]<=2;
			data[82][11:8]<=11;data[82][7:5]<=2;data[82][4:0]<=2;
			data[83][11:8]<=13;data[83][7:5]<=2;data[83][4:0]<=2;
			data[84][11:8]<=2;data[84][7:5]<=1;data[84][4:0]<=2;
			data[85][11:8]<=13;data[85][7:5]<=2;data[85][4:0]<=4;
			data[86][11:8]<=4;data[86][7:5]<=1;data[86][4:0]<=4;
			data[87][11:8]<=2;data[87][7:5]<=1;data[87][4:0]<=4;
			data[88][11:8]<=11;data[88][7:5]<=2;data[88][4:0]<=4;
			data[89][11:8]<=9;data[89][7:5]<=2;data[89][4:0]<=10;
			data[90][11:8]<=0;data[90][7:5]<=2;data[90][4:0]<=2;
			data[91][11:8]<=6;data[91][7:5]<=1;data[91][4:0]<=3;
			data[92][11:8]<=4;data[92][7:5]<=1;data[92][4:0]<=1;
			data[93][11:8]<=2;data[93][7:5]<=1;data[93][4:0]<=8;
			data[94][11:8]<=9;data[94][7:5]<=2;data[94][4:0]<=4;
			data[95][11:8]<=6;data[95][7:5]<=2;data[95][4:0]<=2;
			data[96][11:8]<=11;data[96][7:5]<=2;data[96][4:0]<=8;
			data[97][11:8]<=7;data[97][7:5]<=2;data[97][4:0]<=2;
			data[98][11:8]<=0;data[98][7:5]<=2;data[98][4:0]<=2;
			data[99][11:8]<=4;data[99][7:5]<=1;data[99][4:0]<=2;
			data[100][11:8]<=2;data[100][7:5]<=1;data[100][4:0]<=1;
			data[101][11:8]<=13;data[101][7:5]<=2;data[101][4:0]<=8;
			data[102][11:8]<=11;data[102][7:5]<=2;data[102][4:0]<=4;
			data[103][11:8]<=9;data[103][7:5]<=2;data[103][4:0]<=4;
			data[104][11:8]<=9;data[104][7:5]<=2;data[104][4:0]<=10;
			data[105][11:8]<=0;data[105][7:5]<=2;data[105][4:0]<=2;
			data[106][11:8]<=9;data[106][7:5]<=2;data[106][4:0]<=4;
			data[107][11:8]<=6;data[107][7:5]<=1;data[107][4:0]<=8;
			data[108][11:8]<=4;data[108][7:5]<=1;data[108][4:0]<=4;
			data[109][11:8]<=9;data[109][7:5]<=2;data[109][4:0]<=4;
			data[110][11:8]<=2;data[110][7:5]<=1;data[110][4:0]<=4;
			data[111][11:8]<=0;data[111][7:5]<=2;data[111][4:0]<=4;
			data[112][11:8]<=13;data[112][7:5]<=2;data[112][4:0]<=6;
			data[113][11:8]<=13;data[113][7:5]<=2;data[113][4:0]<=2;
			data[114][11:8]<=11;data[114][7:5]<=2;data[114][4:0]<=6;
			data[115][11:8]<=10;data[115][7:5]<=2;data[115][4:0]<=2;
			data[116][11:8]<=11;data[116][7:5]<=2;data[116][4:0]<=4;
			data[117][11:8]<=4;data[117][7:5]<=1;data[117][4:0]<=4;
			data[118][11:8]<=4;data[118][7:5]<=1;data[118][4:0]<=10;
			data[119][11:8]<=0;data[119][7:5]<=2;data[119][4:0]<=0;
			data[120][11:8]<=6;data[120][7:5]<=1;data[120][4:0]<=2;
			data[121][11:8]<=4;data[121][7:5]<=1;data[121][4:0]<=1;
			data[122][11:8]<=2;data[122][7:5]<=1;data[122][4:0]<=8;
			data[123][11:8]<=9;data[123][7:5]<=2;data[123][4:0]<=6;
			data[124][11:8]<=6;data[124][7:5]<=2;data[124][4:0]<=2;
			data[125][11:8]<=11;data[125][7:5]<=2;data[125][4:0]<=8;
			data[126][11:8]<=7;data[126][7:5]<=2;data[126][4:0]<=2;
			data[127][11:8]<=0;data[127][7:5]<=2;data[127][4:0]<=2;
			data[128][11:8]<=4;data[128][7:5]<=2;data[128][4:0]<=3;
			data[129][11:8]<=2;data[129][7:5]<=2;data[129][4:0]<=1;
			data[130][11:8]<=13;data[130][7:5]<=2;data[130][4:0]<=8;
			data[131][11:8]<=11;data[131][7:5]<=2;data[131][4:0]<=4;
			data[132][11:8]<=9;data[132][7:5]<=2;data[132][4:0]<=4;
			data[133][11:8]<=6;data[133][7:5]<=1;data[133][4:0]<=12;
			data[134][11:8]<=6;data[134][7:5]<=1;data[134][4:0]<=4;
			data[135][11:8]<=9;data[135][7:5]<=1;data[135][4:0]<=8;
			data[136][11:8]<=7;data[136][7:5]<=1;data[136][4:0]<=4;
			data[137][11:8]<=6;data[137][7:5]<=1;data[137][4:0]<=4;
			data[138][11:8]<=4;data[138][7:5]<=1;data[138][4:0]<=6;
			data[139][11:8]<=6;data[139][7:5]<=1;data[139][4:0]<=2;
			data[140][11:8]<=7;data[140][7:5]<=1;data[140][4:0]<=4;
			data[141][11:8]<=0;data[141][7:5]<=2;data[141][4:0]<=2;
			data[142][11:8]<=7;data[142][7:5]<=1;data[142][4:0]<=2;
			data[143][11:8]<=6;data[143][7:5]<=1;data[143][4:0]<=6;
			data[144][11:8]<=6;data[144][7:5]<=1;data[144][4:0]<=2;
			data[145][11:8]<=4;data[145][7:5]<=1;data[145][4:0]<=6;
			data[146][11:8]<=4;data[146][7:5]<=1;data[146][4:0]<=2;
			data[147][11:8]<=2;data[147][7:5]<=1;data[147][4:0]<=12;
			data[148][11:8]<=9;data[148][7:5]<=2;data[148][4:0]<=4;
			data[149][11:8]<=2;data[149][7:5]<=1;data[149][4:0]<=12;
		end
		else if(wen_c)
			data[addr_c] <= data_c;
	end
	assign q_a = data[addr_a];
	assign q_b = data[addr_b];
	endmodule
