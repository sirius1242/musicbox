`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/23 11:16:25
// Design Name: 
// Module Name: regfile
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module regfile(
    input clk, 
		input rst_n, 
		input [15:0] addr_a, 
		input [15:0] addr_b, 
		input [15:0] addr_c, 
		input [11:0] data_c, 
		input wen_c,
		input [2:0] sel,
		output wire [11:0] q_a, 
		output wire [11:0] q_b,
		output [2:0] len,
		output [15:0] addr_d
	);
	integer i;
	reg [11:0] data [0:1000];
	wire [15:0] addr [0:3];
	assign len = 3'b011;
	assign addr[0] = 0;
	assign addr[1] = 152;
	assign addr[2] = 317;
	assign addr[3] = 711;
	assign addr_d = addr[sel];
	always@(posedge clk or negedge rst_n)
	begin
		if (~rst_n)
		begin
			data[0][11:8]<=0;data[0][7:5]<=4;data[0][4:0]<=4;
			data[1][11:8]<=0;data[1][7:5]<=4;data[1][4:0]<=4;
			data[2][11:8]<=0;data[2][7:5]<=4;data[2][4:0]<=4;
			data[3][11:8]<=6;data[3][7:5]<=4;data[3][4:0]<=4;
			data[4][11:8]<=9;data[4][7:5]<=4;data[4][4:0]<=6;
			data[5][11:8]<=9;data[5][7:5]<=4;data[5][4:0]<=2;
			data[6][11:8]<=7;data[6][7:5]<=4;data[6][4:0]<=4;
			data[7][11:8]<=6;data[7][7:5]<=4;data[7][4:0]<=4;
			data[8][11:8]<=4;data[8][7:5]<=4;data[8][4:0]<=6;
			data[9][11:8]<=6;data[9][7:5]<=4;data[9][4:0]<=2;
			data[10][11:8]<=7;data[10][7:5]<=4;data[10][4:0]<=6;
			data[11][11:8]<=7;data[11][7:5]<=4;data[11][4:0]<=2;
			data[12][11:8]<=6;data[12][7:5]<=4;data[12][4:0]<=6;
			data[13][11:8]<=6;data[13][7:5]<=4;data[13][4:0]<=2;
			data[14][11:8]<=4;data[14][7:5]<=4;data[14][4:0]<=6;
			data[15][11:8]<=4;data[15][7:5]<=4;data[15][4:0]<=2;
			data[16][11:8]<=2;data[16][7:5]<=4;data[16][4:0]<=12;
			data[17][11:8]<=9;data[17][7:5]<=4;data[17][4:0]<=4;
			data[18][11:8]<=2;data[18][7:5]<=3;data[18][4:0]<=6;
			data[19][11:8]<=13;data[19][7:5]<=4;data[19][4:0]<=2;
			data[20][11:8]<=4;data[20][7:5]<=3;data[20][4:0]<=2;
			data[21][11:8]<=2;data[21][7:5]<=3;data[21][4:0]<=2;
			data[22][11:8]<=9;data[22][7:5]<=4;data[22][4:0]<=2;
			data[23][11:8]<=6;data[23][7:5]<=4;data[23][4:0]<=2;
			data[24][11:8]<=11;data[24][7:5]<=4;data[24][4:0]<=8;
			data[25][11:8]<=7;data[25][7:5]<=4;data[25][4:0]<=4;
			data[26][11:8]<=0;data[26][7:5]<=4;data[26][4:0]<=2;
			data[27][11:8]<=11;data[27][7:5]<=4;data[27][4:0]<=2;
			data[28][11:8]<=4;data[28][7:5]<=3;data[28][4:0]<=6;
			data[29][11:8]<=2;data[29][7:5]<=4;data[29][4:0]<=4;
			data[30][11:8]<=13;data[30][7:5]<=4;data[30][4:0]<=2;
			data[31][11:8]<=11;data[31][7:5]<=4;data[31][4:0]<=2;
			data[32][11:8]<=9;data[32][7:5]<=4;data[32][4:0]<=2;
			data[33][11:8]<=7;data[33][7:5]<=4;data[33][4:0]<=2;
			data[34][11:8]<=6;data[34][7:5]<=4;data[34][4:0]<=12;
			data[35][11:8]<=9;data[35][7:5]<=4;data[35][4:0]<=2;
			data[36][11:8]<=2;data[36][7:5]<=3;data[36][4:0]<=6;
			data[37][11:8]<=13;data[37][7:5]<=4;data[37][4:0]<=2;
			data[38][11:8]<=4;data[38][7:5]<=3;data[38][4:0]<=2;
			data[39][11:8]<=2;data[39][7:5]<=3;data[39][4:0]<=2;
			data[40][11:8]<=9;data[40][7:5]<=4;data[40][4:0]<=2;
			data[41][11:8]<=6;data[41][7:5]<=4;data[41][4:0]<=2;
			data[42][11:8]<=11;data[42][7:5]<=4;data[42][4:0]<=8;
			data[43][11:8]<=7;data[43][7:5]<=4;data[43][4:0]<=2;
			data[44][11:8]<=11;data[44][7:5]<=4;data[44][4:0]<=2;
			data[45][11:8]<=4;data[45][7:5]<=3;data[45][4:0]<=2;
			data[46][11:8]<=2;data[46][7:5]<=3;data[46][4:0]<=2;
			data[47][11:8]<=13;data[47][7:5]<=4;data[47][4:0]<=4;
			data[48][11:8]<=4;data[48][7:5]<=3;data[48][4:0]<=4;
			data[49][11:8]<=7;data[49][7:5]<=3;data[49][4:0]<=4;
			data[50][11:8]<=13;data[50][7:5]<=4;data[50][4:0]<=4;
			data[51][11:8]<=2;data[51][7:5]<=3;data[51][4:0]<=8;
			data[52][11:8]<=2;data[52][7:5]<=3;data[52][4:0]<=2;
			data[53][11:8]<=0;data[53][7:5]<=4;data[53][4:0]<=2;
			data[54][11:8]<=6;data[54][7:5]<=3;data[54][4:0]<=2;
			data[55][11:8]<=4;data[55][7:5]<=3;data[55][4:0]<=2;
			data[56][11:8]<=13;data[56][7:5]<=4;data[56][4:0]<=8;
			data[57][11:8]<=11;data[57][7:5]<=4;data[57][4:0]<=2;
			data[58][11:8]<=13;data[58][7:5]<=4;data[58][4:0]<=2;
			data[59][11:8]<=2;data[59][7:5]<=3;data[59][4:0]<=2;
			data[60][11:8]<=11;data[60][7:5]<=4;data[60][4:0]<=2;
			data[61][11:8]<=13;data[61][7:5]<=4;data[61][4:0]<=8;
			data[62][11:8]<=9;data[62][7:5]<=4;data[62][4:0]<=2;
			data[63][11:8]<=9;data[63][7:5]<=4;data[63][4:0]<=2;
			data[64][11:8]<=8;data[64][7:5]<=4;data[64][4:0]<=2;
			data[65][11:8]<=9;data[65][7:5]<=4;data[65][4:0]<=2;
			data[66][11:8]<=11;data[66][7:5]<=4;data[66][4:0]<=6;
			data[67][11:8]<=11;data[67][7:5]<=4;data[67][4:0]<=2;
			data[68][11:8]<=4;data[68][7:5]<=3;data[68][4:0]<=4;
			data[69][11:8]<=2;data[69][7:5]<=3;data[69][4:0]<=2;
			data[70][11:8]<=13;data[70][7:5]<=4;data[70][4:0]<=8;
			data[71][11:8]<=13;data[71][7:5]<=4;data[71][4:0]<=2;
			data[72][11:8]<=0;data[72][7:5]<=4;data[72][4:0]<=2;
			data[73][11:8]<=4;data[73][7:5]<=3;data[73][4:0]<=4;
			data[74][11:8]<=4;data[74][7:5]<=3;data[74][4:0]<=6;
			data[75][11:8]<=13;data[75][7:5]<=4;data[75][4:0]<=2;
			data[76][11:8]<=9;data[76][7:5]<=4;data[76][4:0]<=2;
			data[77][11:8]<=9;data[77][7:5]<=4;data[77][4:0]<=2;
			data[78][11:8]<=8;data[78][7:5]<=4;data[78][4:0]<=2;
			data[79][11:8]<=9;data[79][7:5]<=4;data[79][4:0]<=2;
			data[80][11:8]<=6;data[80][7:5]<=3;data[80][4:0]<=8;
			data[81][11:8]<=2;data[81][7:5]<=3;data[81][4:0]<=2;
			data[82][11:8]<=11;data[82][7:5]<=4;data[82][4:0]<=2;
			data[83][11:8]<=13;data[83][7:5]<=4;data[83][4:0]<=2;
			data[84][11:8]<=2;data[84][7:5]<=3;data[84][4:0]<=2;
			data[85][11:8]<=13;data[85][7:5]<=4;data[85][4:0]<=4;
			data[86][11:8]<=4;data[86][7:5]<=3;data[86][4:0]<=4;
			data[87][11:8]<=2;data[87][7:5]<=3;data[87][4:0]<=4;
			data[88][11:8]<=11;data[88][7:5]<=4;data[88][4:0]<=4;
			data[89][11:8]<=9;data[89][7:5]<=4;data[89][4:0]<=10;
			data[90][11:8]<=0;data[90][7:5]<=4;data[90][4:0]<=2;
			data[91][11:8]<=6;data[91][7:5]<=3;data[91][4:0]<=3;
			data[92][11:8]<=4;data[92][7:5]<=3;data[92][4:0]<=1;
			data[93][11:8]<=2;data[93][7:5]<=3;data[93][4:0]<=8;
			data[94][11:8]<=9;data[94][7:5]<=4;data[94][4:0]<=4;
			data[95][11:8]<=6;data[95][7:5]<=4;data[95][4:0]<=2;
			data[96][11:8]<=11;data[96][7:5]<=4;data[96][4:0]<=8;
			data[97][11:8]<=7;data[97][7:5]<=4;data[97][4:0]<=2;
			data[98][11:8]<=0;data[98][7:5]<=4;data[98][4:0]<=2;
			data[99][11:8]<=4;data[99][7:5]<=3;data[99][4:0]<=2;
			data[100][11:8]<=2;data[100][7:5]<=3;data[100][4:0]<=1;
			data[101][11:8]<=13;data[101][7:5]<=4;data[101][4:0]<=8;
			data[102][11:8]<=11;data[102][7:5]<=4;data[102][4:0]<=4;
			data[103][11:8]<=9;data[103][7:5]<=4;data[103][4:0]<=4;
			data[104][11:8]<=9;data[104][7:5]<=4;data[104][4:0]<=10;
			data[105][11:8]<=0;data[105][7:5]<=4;data[105][4:0]<=2;
			data[106][11:8]<=9;data[106][7:5]<=4;data[106][4:0]<=4;
			data[107][11:8]<=6;data[107][7:5]<=3;data[107][4:0]<=8;
			data[108][11:8]<=4;data[108][7:5]<=3;data[108][4:0]<=4;
			data[109][11:8]<=9;data[109][7:5]<=4;data[109][4:0]<=4;
			data[110][11:8]<=2;data[110][7:5]<=3;data[110][4:0]<=4;
			data[111][11:8]<=0;data[111][7:5]<=4;data[111][4:0]<=4;
			data[112][11:8]<=13;data[112][7:5]<=4;data[112][4:0]<=6;
			data[113][11:8]<=13;data[113][7:5]<=4;data[113][4:0]<=2;
			data[114][11:8]<=11;data[114][7:5]<=4;data[114][4:0]<=6;
			data[115][11:8]<=10;data[115][7:5]<=4;data[115][4:0]<=2;
			data[116][11:8]<=11;data[116][7:5]<=4;data[116][4:0]<=4;
			data[117][11:8]<=4;data[117][7:5]<=3;data[117][4:0]<=4;
			data[118][11:8]<=4;data[118][7:5]<=3;data[118][4:0]<=10;
			data[119][11:8]<=0;data[119][7:5]<=4;data[119][4:0]<=2;
			data[120][11:8]<=6;data[120][7:5]<=3;data[120][4:0]<=2;
			data[121][11:8]<=4;data[121][7:5]<=3;data[121][4:0]<=1;
			data[122][11:8]<=2;data[122][7:5]<=3;data[122][4:0]<=8;
			data[123][11:8]<=9;data[123][7:5]<=4;data[123][4:0]<=6;
			data[124][11:8]<=6;data[124][7:5]<=4;data[124][4:0]<=2;
			data[125][11:8]<=11;data[125][7:5]<=4;data[125][4:0]<=8;
			data[126][11:8]<=7;data[126][7:5]<=4;data[126][4:0]<=2;
			data[127][11:8]<=0;data[127][7:5]<=4;data[127][4:0]<=2;
			data[128][11:8]<=4;data[128][7:5]<=4;data[128][4:0]<=3;
			data[129][11:8]<=2;data[129][7:5]<=4;data[129][4:0]<=1;
			data[130][11:8]<=13;data[130][7:5]<=4;data[130][4:0]<=8;
			data[131][11:8]<=11;data[131][7:5]<=4;data[131][4:0]<=4;
			data[132][11:8]<=9;data[132][7:5]<=4;data[132][4:0]<=4;
			data[133][11:8]<=6;data[133][7:5]<=3;data[133][4:0]<=12;
			data[134][11:8]<=6;data[134][7:5]<=3;data[134][4:0]<=4;
			data[135][11:8]<=9;data[135][7:5]<=3;data[135][4:0]<=8;
			data[136][11:8]<=7;data[136][7:5]<=3;data[136][4:0]<=4;
			data[137][11:8]<=6;data[137][7:5]<=3;data[137][4:0]<=4;
			data[138][11:8]<=4;data[138][7:5]<=3;data[138][4:0]<=6;
			data[139][11:8]<=6;data[139][7:5]<=3;data[139][4:0]<=2;
			data[140][11:8]<=7;data[140][7:5]<=3;data[140][4:0]<=4;
			data[141][11:8]<=0;data[141][7:5]<=4;data[141][4:0]<=2;
			data[142][11:8]<=7;data[142][7:5]<=3;data[142][4:0]<=2;
			data[143][11:8]<=6;data[143][7:5]<=3;data[143][4:0]<=6;
			data[144][11:8]<=6;data[144][7:5]<=3;data[144][4:0]<=2;
			data[145][11:8]<=4;data[145][7:5]<=3;data[145][4:0]<=6;
			data[146][11:8]<=4;data[146][7:5]<=3;data[146][4:0]<=2;
			data[147][11:8]<=2;data[147][7:5]<=3;data[147][4:0]<=12;
			data[148][11:8]<=9;data[148][7:5]<=4;data[148][4:0]<=4;
			data[149][11:8]<=2;data[149][7:5]<=3;data[149][4:0]<=12;

			data[152][11:8]<=0;data[152][7:5]<=4;data[152][4:0]<=4;
			data[153][11:8]<=0;data[153][7:5]<=4;data[153][4:0]<=4;
			data[154][11:8]<=0;data[154][7:5]<=4;data[154][4:0]<=4;
			data[155][11:8]<=0;data[155][7:5]<=4;data[155][4:0]<=4;
			data[156][11:8]<=0;data[156][7:5]<=4;data[156][4:0]<=2;
			data[157][11:8]<=6;data[157][7:5]<=4;data[157][4:0]<=2;
			data[158][11:8]<=6;data[158][7:5]<=4;data[158][4:0]<=2;
			data[159][11:8]<=6;data[159][7:5]<=4;data[159][4:0]<=2;
			data[160][11:8]<=6;data[160][7:5]<=4;data[160][4:0]<=2;
			data[161][11:8]<=4;data[161][7:5]<=4;data[161][4:0]<=2;
			data[162][11:8]<=6;data[162][7:5]<=4;data[162][4:0]<=2;
			data[163][11:8]<=11;data[163][7:5]<=4;data[163][4:0]<=2;
			data[164][11:8]<=6;data[164][7:5]<=4;data[164][4:0]<=2;
			data[165][11:8]<=4;data[165][7:5]<=4;data[165][4:0]<=1;
			data[166][11:8]<=4;data[166][7:5]<=4;data[166][4:0]<=5;
			data[167][11:8]<=0;data[167][7:5]<=4;data[167][4:0]<=4;
			data[168][11:8]<=0;data[168][7:5]<=4;data[168][4:0]<=4;
			data[169][11:8]<=0;data[169][7:5]<=4;data[169][4:0]<=2;
			data[170][11:8]<=4;data[170][7:5]<=4;data[170][4:0]<=2;
			data[171][11:8]<=4;data[171][7:5]<=4;data[171][4:0]<=2;
			data[172][11:8]<=4;data[172][7:5]<=4;data[172][4:0]<=2;
			data[173][11:8]<=4;data[173][7:5]<=4;data[173][4:0]<=2;
			data[174][11:8]<=2;data[174][7:5]<=4;data[174][4:0]<=2;
			data[175][11:8]<=4;data[175][7:5]<=4;data[175][4:0]<=2;
			data[176][11:8]<=9;data[176][7:5]<=4;data[176][4:0]<=2;
			data[177][11:8]<=4;data[177][7:5]<=4;data[177][4:0]<=2;
			data[178][11:8]<=2;data[178][7:5]<=4;data[178][4:0]<=2;
			data[179][11:8]<=13;data[179][7:5]<=5;data[179][4:0]<=2;
			data[180][11:8]<=2;data[180][7:5]<=4;data[180][4:0]<=6;
			data[181][11:8]<=0;data[181][7:5]<=4;data[181][4:0]<=2;
			data[182][11:8]<=11;data[182][7:5]<=5;data[182][4:0]<=1;
			data[183][11:8]<=13;data[183][7:5]<=5;data[183][4:0]<=1;
			data[184][11:8]<=2;data[184][7:5]<=4;data[184][4:0]<=2;
			data[185][11:8]<=2;data[185][7:5]<=4;data[185][4:0]<=2;
			data[186][11:8]<=2;data[186][7:5]<=4;data[186][4:0]<=2;
			data[187][11:8]<=2;data[187][7:5]<=4;data[187][4:0]<=2;
			data[188][11:8]<=2;data[188][7:5]<=4;data[188][4:0]<=4;
			data[189][11:8]<=0;data[189][7:5]<=4;data[189][4:0]<=2;
			data[190][11:8]<=11;data[190][7:5]<=5;data[190][4:0]<=1;
			data[191][11:8]<=13;data[191][7:5]<=5;data[191][4:0]<=1;
			data[192][11:8]<=2;data[192][7:5]<=4;data[192][4:0]<=2;
			data[193][11:8]<=2;data[193][7:5]<=4;data[193][4:0]<=2;
			data[194][11:8]<=2;data[194][7:5]<=4;data[194][4:0]<=2;
			data[195][11:8]<=2;data[195][7:5]<=4;data[195][4:0]<=2;
			data[196][11:8]<=13;data[196][7:5]<=5;data[196][4:0]<=2;
			data[197][11:8]<=2;data[197][7:5]<=4;data[197][4:0]<=2;
			data[198][11:8]<=0;data[198][7:5]<=4;data[198][4:0]<=2;
			data[199][11:8]<=11;data[199][7:5]<=5;data[199][4:0]<=1;
			data[200][11:8]<=13;data[200][7:5]<=5;data[200][4:0]<=1;
			data[201][11:8]<=2;data[201][7:5]<=4;data[201][4:0]<=2;
			data[202][11:8]<=2;data[202][7:5]<=4;data[202][4:0]<=2;
			data[203][11:8]<=2;data[203][7:5]<=4;data[203][4:0]<=2;
			data[204][11:8]<=2;data[204][7:5]<=4;data[204][4:0]<=2;
			data[205][11:8]<=2;data[205][7:5]<=4;data[205][4:0]<=2;
			data[206][11:8]<=9;data[206][7:5]<=4;data[206][4:0]<=4;
			data[207][11:8]<=2;data[207][7:5]<=4;data[207][4:0]<=2;
			data[208][11:8]<=4;data[208][7:5]<=4;data[208][4:0]<=8;
			data[209][11:8]<=6;data[209][7:5]<=4;data[209][4:0]<=4;
			data[210][11:8]<=7;data[210][7:5]<=4;data[210][4:0]<=4;
			data[211][11:8]<=9;data[211][7:5]<=4;data[211][4:0]<=2;
			data[212][11:8]<=9;data[212][7:5]<=4;data[212][4:0]<=4;
			data[213][11:8]<=9;data[213][7:5]<=4;data[213][4:0]<=2;
			data[214][11:8]<=9;data[214][7:5]<=4;data[214][4:0]<=2;
			data[215][11:8]<=7;data[215][7:5]<=4;data[215][4:0]<=2;
			data[216][11:8]<=6;data[216][7:5]<=4;data[216][4:0]<=2;
			data[217][11:8]<=4;data[217][7:5]<=4;data[217][4:0]<=2;
			data[218][11:8]<=4;data[218][7:5]<=4;data[218][4:0]<=2;
			data[219][11:8]<=6;data[219][7:5]<=4;data[219][4:0]<=1;
			data[220][11:8]<=2;data[220][7:5]<=4;data[220][4:0]<=5;
			data[221][11:8]<=0;data[221][7:5]<=4;data[221][4:0]<=4;
			data[222][11:8]<=6;data[222][7:5]<=4;data[222][4:0]<=2;
			data[223][11:8]<=7;data[223][7:5]<=4;data[223][4:0]<=2;
			data[224][11:8]<=9;data[224][7:5]<=4;data[224][4:0]<=2;
			data[225][11:8]<=9;data[225][7:5]<=6;data[225][4:0]<=4;
			data[226][11:8]<=9;data[226][7:5]<=4;data[226][4:0]<=2;
			data[227][11:8]<=9;data[227][7:5]<=4;data[227][4:0]<=2;
			data[228][11:8]<=7;data[228][7:5]<=4;data[228][4:0]<=2;
			data[229][11:8]<=6;data[229][7:5]<=4;data[229][4:0]<=2;
			data[230][11:8]<=4;data[230][7:5]<=4;data[230][4:0]<=2;
			data[231][11:8]<=4;data[231][7:5]<=4;data[231][4:0]<=2;
			data[232][11:8]<=6;data[232][7:5]<=4;data[232][4:0]<=10;
			data[233][11:8]<=2;data[233][7:5]<=4;data[233][4:0]<=2;
			data[234][11:8]<=4;data[234][7:5]<=4;data[234][4:0]<=2;
			data[235][11:8]<=6;data[235][7:5]<=4;data[235][4:0]<=6;
			data[236][11:8]<=11;data[236][7:5]<=5;data[236][4:0]<=2;
			data[237][11:8]<=2;data[237][7:5]<=4;data[237][4:0]<=2;
			data[238][11:8]<=13;data[238][7:5]<=5;data[238][4:0]<=2;
			data[239][11:8]<=2;data[239][7:5]<=4;data[239][4:0]<=2;
			data[240][11:8]<=6;data[240][7:5]<=4;data[240][4:0]<=8;
			data[241][11:8]<=4;data[241][7:5]<=4;data[241][4:0]<=4;
			data[242][11:8]<=11;data[242][7:5]<=4;data[242][4:0]<=2;
			data[243][11:8]<=13;data[243][7:5]<=4;data[243][4:0]<=2;
			data[244][11:8]<=2;data[244][7:5]<=3;data[244][4:0]<=2;
			data[245][11:8]<=2;data[245][7:5]<=3;data[245][4:0]<=2;
			data[246][11:8]<=4;data[246][7:5]<=3;data[246][4:0]<=2;
			data[247][11:8]<=2;data[247][7:5]<=3;data[247][4:0]<=2;
			data[248][11:8]<=13;data[248][7:5]<=4;data[248][4:0]<=4;
			data[249][11:8]<=6;data[249][7:5]<=4;data[249][4:0]<=2;
			data[250][11:8]<=9;data[250][7:5]<=4;data[250][4:0]<=2;
			data[251][11:8]<=11;data[251][7:5]<=4;data[251][4:0]<=2;
			data[252][11:8]<=11;data[252][7:5]<=4;data[252][4:0]<=2;
			data[253][11:8]<=9;data[253][7:5]<=4;data[253][4:0]<=2;
			data[254][11:8]<=7;data[254][7:5]<=4;data[254][4:0]<=2;
			data[255][11:8]<=9;data[255][7:5]<=4;data[255][4:0]<=6;
			data[256][11:8]<=9;data[256][7:5]<=4;data[256][4:0]<=2;
			data[257][11:8]<=9;data[257][7:5]<=4;data[257][4:0]<=2;
			data[258][11:8]<=7;data[258][7:5]<=4;data[258][4:0]<=2;
			data[259][11:8]<=7;data[259][7:5]<=4;data[259][4:0]<=2;
			data[260][11:8]<=5;data[260][7:5]<=4;data[260][4:0]<=2;
			data[261][11:8]<=7;data[261][7:5]<=4;data[261][4:0]<=4;
			data[262][11:8]<=2;data[262][7:5]<=4;data[262][4:0]<=2;
			data[263][11:8]<=7;data[263][7:5]<=4;data[263][4:0]<=2;
			data[264][11:8]<=9;data[264][7:5]<=4;data[264][4:0]<=6;
			data[265][11:8]<=10;data[265][7:5]<=4;data[265][4:0]<=2;
			data[266][11:8]<=9;data[266][7:5]<=4;data[266][4:0]<=4;
			data[267][11:8]<=11;data[267][7:5]<=4;data[267][4:0]<=2;
			data[268][11:8]<=13;data[268][7:5]<=4;data[268][4:0]<=2;
			data[269][11:8]<=2;data[269][7:5]<=3;data[269][4:0]<=2;
			data[270][11:8]<=2;data[270][7:5]<=3;data[270][4:0]<=2;
			data[271][11:8]<=4;data[271][7:5]<=3;data[271][4:0]<=2;
			data[272][11:8]<=2;data[272][7:5]<=3;data[272][4:0]<=2;
			data[273][11:8]<=13;data[273][7:5]<=4;data[273][4:0]<=4;
			data[274][11:8]<=6;data[274][7:5]<=4;data[274][4:0]<=2;
			data[275][11:8]<=9;data[275][7:5]<=4;data[275][4:0]<=2;
			data[276][11:8]<=11;data[276][7:5]<=4;data[276][4:0]<=2;
			data[277][11:8]<=11;data[277][7:5]<=4;data[277][4:0]<=2;
			data[278][11:8]<=9;data[278][7:5]<=4;data[278][4:0]<=2;
			data[279][11:8]<=7;data[279][7:5]<=4;data[279][4:0]<=2;
			data[280][11:8]<=9;data[280][7:5]<=4;data[280][4:0]<=6;
			data[281][11:8]<=9;data[281][7:5]<=4;data[281][4:0]<=2;
			data[282][11:8]<=9;data[282][7:5]<=4;data[282][4:0]<=2;
			data[283][11:8]<=7;data[283][7:5]<=4;data[283][4:0]<=2;
			data[284][11:8]<=7;data[284][7:5]<=4;data[284][4:0]<=2;
			data[285][11:8]<=5;data[285][7:5]<=4;data[285][4:0]<=2;
			data[286][11:8]<=7;data[286][7:5]<=4;data[286][4:0]<=4;
			data[287][11:8]<=9;data[287][7:5]<=4;data[287][4:0]<=2;
			data[288][11:8]<=10;data[288][7:5]<=4;data[288][4:0]<=2;
			data[289][11:8]<=12;data[289][7:5]<=4;data[289][4:0]<=2;
			data[290][11:8]<=10;data[290][7:5]<=4;data[290][4:0]<=2;
			data[291][11:8]<=10;data[291][7:5]<=4;data[291][4:0]<=2;
			data[292][11:8]<=9;data[292][7:5]<=4;data[292][4:0]<=2;
			data[293][11:8]<=9;data[293][7:5]<=4;data[293][4:0]<=2;
			data[294][11:8]<=9;data[294][7:5]<=4;data[294][4:0]<=2;
			data[295][11:8]<=10;data[295][7:5]<=4;data[295][4:0]<=2;
			data[296][11:8]<=13;data[296][7:5]<=4;data[296][4:0]<=2;
			data[297][11:8]<=2;data[297][7:5]<=3;data[297][4:0]<=12;
			data[298][11:8]<=10;data[298][7:5]<=4;data[298][4:0]<=2;
			data[299][11:8]<=12;data[299][7:5]<=4;data[299][4:0]<=2;
			data[300][11:8]<=2;data[300][7:5]<=3;data[300][4:0]<=8;
			data[301][11:8]<=0;data[301][7:5]<=4;data[301][4:0]<=2;
			data[302][11:8]<=2;data[302][7:5]<=3;data[302][4:0]<=2;
			data[303][11:8]<=13;data[303][7:5]<=4;data[303][4:0]<=2;
			data[304][11:8]<=2;data[304][7:5]<=3;data[304][4:0]<=2;
			data[305][11:8]<=4;data[305][7:5]<=3;data[305][4:0]<=8;
			data[306][11:8]<=0;data[306][7:5]<=4;data[306][4:0]<=2;
			data[307][11:8]<=9;data[307][7:5]<=4;data[307][4:0]<=2;
			data[308][11:8]<=2;data[308][7:5]<=3;data[308][4:0]<=2;
			data[309][11:8]<=13;data[309][7:5]<=4;data[309][4:0]<=2;
			data[310][11:8]<=2;data[310][7:5]<=3;data[310][4:0]<=16;
			data[311][11:8]<=0;data[311][7:5]<=4;data[311][4:0]<=16;
			data[312][11:8]<=0;data[312][7:5]<=4;data[312][4:0]<=16;
			data[313][11:8]<=0;data[313][7:5]<=4;data[313][4:0]<=16;

			data[317][11:8]<=6;data[317][7:5]<=3;data[317][4:0]<=8;
			data[318][11:8]<=4;data[318][7:5]<=3;data[318][4:0]<=3;
			data[319][11:8]<=2;data[319][7:5]<=3;data[319][4:0]<=8;
			data[320][11:8]<=13;data[320][7:5]<=4;data[320][4:0]<=8;
			data[321][11:8]<=11;data[321][7:5]<=4;data[321][4:0]<=8;
			data[322][11:8]<=9;data[322][7:5]<=4;data[322][4:0]<=8;
			data[323][11:8]<=11;data[323][7:5]<=4;data[323][4:0]<=8;
			data[324][11:8]<=13;data[324][7:5]<=4;data[324][4:0]<=8;
			data[325][11:8]<=2;data[325][7:5]<=3;data[325][4:0]<=8;
			data[326][11:8]<=13;data[326][7:5]<=4;data[326][4:0]<=8;
			data[327][11:8]<=11;data[327][7:5]<=4;data[327][4:0]<=8;
			data[328][11:8]<=9;data[328][7:5]<=4;data[328][4:0]<=8;
			data[329][11:8]<=7;data[329][7:5]<=4;data[329][4:0]<=8;
			data[330][11:8]<=6;data[330][7:5]<=4;data[330][4:0]<=8;
			data[331][11:8]<=7;data[331][7:5]<=4;data[331][4:0]<=8;
			data[332][11:8]<=4;data[332][7:5]<=4;data[332][4:0]<=8;
			data[333][11:8]<=2;data[333][7:5]<=3;data[333][4:0]<=2;
			data[334][11:8]<=13;data[334][7:5]<=4;data[334][4:0]<=2;
			data[335][11:8]<=2;data[335][7:5]<=3;data[335][4:0]<=2;
			data[336][11:8]<=2;data[336][7:5]<=4;data[336][4:0]<=2;
			data[337][11:8]<=13;data[337][7:5]<=5;data[337][4:0]<=2;
			data[338][11:8]<=9;data[338][7:5]<=4;data[338][4:0]<=2;
			data[339][11:8]<=4;data[339][7:5]<=4;data[339][4:0]<=2;
			data[340][11:8]<=6;data[340][7:5]<=4;data[340][4:0]<=2;
			data[341][11:8]<=2;data[341][7:5]<=4;data[341][4:0]<=2;
			data[342][11:8]<=2;data[342][7:5]<=3;data[342][4:0]<=2;
			data[343][11:8]<=13;data[343][7:5]<=4;data[343][4:0]<=2;
			data[344][11:8]<=11;data[344][7:5]<=4;data[344][4:0]<=2;
			data[345][11:8]<=13;data[345][7:5]<=4;data[345][4:0]<=2;
			data[346][11:8]<=6;data[346][7:5]<=3;data[346][4:0]<=2;
			data[347][11:8]<=9;data[347][7:5]<=3;data[347][4:0]<=2;
			data[348][11:8]<=11;data[348][7:5]<=3;data[348][4:0]<=2;
			data[349][11:8]<=7;data[349][7:5]<=3;data[349][4:0]<=2;
			data[350][11:8]<=6;data[350][7:5]<=3;data[350][4:0]<=2;
			data[351][11:8]<=4;data[351][7:5]<=3;data[351][4:0]<=2;
			data[352][11:8]<=7;data[352][7:5]<=3;data[352][4:0]<=2;
			data[353][11:8]<=7;data[353][7:5]<=3;data[353][4:0]<=2;
			data[354][11:8]<=6;data[354][7:5]<=3;data[354][4:0]<=2;
			data[355][11:8]<=2;data[355][7:5]<=3;data[355][4:0]<=2;
			data[356][11:8]<=13;data[356][7:5]<=4;data[356][4:0]<=2;
			data[357][11:8]<=11;data[357][7:5]<=4;data[357][4:0]<=2;
			data[358][11:8]<=9;data[358][7:5]<=4;data[358][4:0]<=2;
			data[359][11:8]<=7;data[359][7:5]<=4;data[359][4:0]<=2;
			data[360][11:8]<=6;data[360][7:5]<=4;data[360][4:0]<=2;
			data[361][11:8]<=4;data[361][7:5]<=4;data[361][4:0]<=2;
			data[362][11:8]<=7;data[362][7:5]<=4;data[362][4:0]<=2;
			data[363][11:8]<=6;data[363][7:5]<=4;data[363][4:0]<=2;
			data[364][11:8]<=4;data[364][7:5]<=4;data[364][4:0]<=2;
			data[365][11:8]<=2;data[365][7:5]<=4;data[365][4:0]<=2;
			data[366][11:8]<=4;data[366][7:5]<=4;data[366][4:0]<=2;
			data[367][11:8]<=6;data[367][7:5]<=4;data[367][4:0]<=2;
			data[368][11:8]<=7;data[368][7:5]<=4;data[368][4:0]<=2;
			data[369][11:8]<=9;data[369][7:5]<=4;data[369][4:0]<=2;
			data[370][11:8]<=4;data[370][7:5]<=4;data[370][4:0]<=2;
			data[371][11:8]<=9;data[371][7:5]<=4;data[371][4:0]<=2;
			data[372][11:8]<=7;data[372][7:5]<=4;data[372][4:0]<=2;
			data[373][11:8]<=6;data[373][7:5]<=4;data[373][4:0]<=2;
			data[374][11:8]<=11;data[374][7:5]<=4;data[374][4:0]<=2;
			data[375][11:8]<=9;data[375][7:5]<=4;data[375][4:0]<=2;
			data[376][11:8]<=7;data[376][7:5]<=4;data[376][4:0]<=2;
			data[377][11:8]<=9;data[377][7:5]<=4;data[377][4:0]<=2;
			data[378][11:8]<=7;data[378][7:5]<=4;data[378][4:0]<=2;
			data[379][11:8]<=6;data[379][7:5]<=4;data[379][4:0]<=2;
			data[380][11:8]<=4;data[380][7:5]<=4;data[380][4:0]<=2;
			data[381][11:8]<=2;data[381][7:5]<=4;data[381][4:0]<=2;
			data[382][11:8]<=11;data[382][7:5]<=5;data[382][4:0]<=2;
			data[383][11:8]<=11;data[383][7:5]<=4;data[383][4:0]<=2;
			data[384][11:8]<=13;data[384][7:5]<=4;data[384][4:0]<=2;
			data[385][11:8]<=2;data[385][7:5]<=3;data[385][4:0]<=2;
			data[386][11:8]<=13;data[386][7:5]<=4;data[386][4:0]<=2;
			data[387][11:8]<=11;data[387][7:5]<=4;data[387][4:0]<=2;
			data[388][11:8]<=9;data[388][7:5]<=4;data[388][4:0]<=2;
			data[389][11:8]<=7;data[389][7:5]<=4;data[389][4:0]<=2;
			data[390][11:8]<=6;data[390][7:5]<=4;data[390][4:0]<=2;
			data[391][11:8]<=4;data[391][7:5]<=4;data[391][4:0]<=2;
			data[392][11:8]<=11;data[392][7:5]<=4;data[392][4:0]<=2;
			data[393][11:8]<=9;data[393][7:5]<=4;data[393][4:0]<=2;
			data[394][11:8]<=11;data[394][7:5]<=4;data[394][4:0]<=2;
			data[395][11:8]<=9;data[395][7:5]<=4;data[395][4:0]<=2;
			data[396][11:8]<=7;data[396][7:5]<=4;data[396][4:0]<=2;
			data[397][11:8]<=6;data[397][7:5]<=4;data[397][4:0]<=4;
			data[398][11:8]<=6;data[398][7:5]<=3;data[398][4:0]<=4;
			data[399][11:8]<=4;data[399][7:5]<=3;data[399][4:0]<=8;
			data[400][11:8]<=2;data[400][7:5]<=3;data[400][4:0]<=8;
			data[401][11:8]<=4;data[401][7:5]<=3;data[401][4:0]<=8;
			data[402][11:8]<=2;data[402][7:5]<=3;data[402][4:0]<=4;
			data[403][11:8]<=6;data[403][7:5]<=3;data[403][4:0]<=4;
			data[404][11:8]<=4;data[404][7:5]<=3;data[404][4:0]<=4;
			data[405][11:8]<=7;data[405][7:5]<=3;data[405][4:0]<=4;
			data[406][11:8]<=9;data[406][7:5]<=3;data[406][4:0]<=2;
			data[407][11:8]<=6;data[407][7:5]<=3;data[407][4:0]<=1;
			data[408][11:8]<=7;data[408][7:5]<=3;data[408][4:0]<=1;
			data[409][11:8]<=9;data[409][7:5]<=3;data[409][4:0]<=2;
			data[410][11:8]<=6;data[410][7:5]<=3;data[410][4:0]<=1;
			data[411][11:8]<=7;data[411][7:5]<=3;data[411][4:0]<=1;
			data[412][11:8]<=9;data[412][7:5]<=3;data[412][4:0]<=1;
			data[413][11:8]<=9;data[413][7:5]<=4;data[413][4:0]<=1;
			data[414][11:8]<=11;data[414][7:5]<=4;data[414][4:0]<=1;
			data[415][11:8]<=13;data[415][7:5]<=4;data[415][4:0]<=1;
			data[416][11:8]<=2;data[416][7:5]<=3;data[416][4:0]<=1;
			data[417][11:8]<=4;data[417][7:5]<=3;data[417][4:0]<=1;
			data[418][11:8]<=6;data[418][7:5]<=3;data[418][4:0]<=1;
			data[419][11:8]<=7;data[419][7:5]<=3;data[419][4:0]<=1;
			data[420][11:8]<=6;data[420][7:5]<=3;data[420][4:0]<=2;
			data[421][11:8]<=2;data[421][7:5]<=3;data[421][4:0]<=1;
			data[422][11:8]<=4;data[422][7:5]<=3;data[422][4:0]<=1;
			data[423][11:8]<=6;data[423][7:5]<=3;data[423][4:0]<=2;
			data[424][11:8]<=6;data[424][7:5]<=4;data[424][4:0]<=1;
			data[425][11:8]<=7;data[425][7:5]<=4;data[425][4:0]<=1;
			data[426][11:8]<=9;data[426][7:5]<=4;data[426][4:0]<=1;
			data[427][11:8]<=11;data[427][7:5]<=4;data[427][4:0]<=1;
			data[428][11:8]<=9;data[428][7:5]<=4;data[428][4:0]<=1;
			data[429][11:8]<=7;data[429][7:5]<=4;data[429][4:0]<=1;
			data[430][11:8]<=9;data[430][7:5]<=4;data[430][4:0]<=1;
			data[431][11:8]<=6;data[431][7:5]<=4;data[431][4:0]<=1;
			data[432][11:8]<=7;data[432][7:5]<=4;data[432][4:0]<=1;
			data[433][11:8]<=9;data[433][7:5]<=4;data[433][4:0]<=1;
			data[434][11:8]<=7;data[434][7:5]<=4;data[434][4:0]<=2;
			data[435][11:8]<=11;data[435][7:5]<=4;data[435][4:0]<=1;
			data[436][11:8]<=9;data[436][7:5]<=4;data[436][4:0]<=1;
			data[437][11:8]<=7;data[437][7:5]<=4;data[437][4:0]<=2;
			data[438][11:8]<=6;data[438][7:5]<=4;data[438][4:0]<=1;
			data[439][11:8]<=4;data[439][7:5]<=4;data[439][4:0]<=1;
			data[440][11:8]<=6;data[440][7:5]<=4;data[440][4:0]<=1;
			data[441][11:8]<=4;data[441][7:5]<=4;data[441][4:0]<=1;
			data[442][11:8]<=2;data[442][7:5]<=4;data[442][4:0]<=1;
			data[443][11:8]<=4;data[443][7:5]<=4;data[443][4:0]<=1;
			data[444][11:8]<=6;data[444][7:5]<=4;data[444][4:0]<=1;
			data[445][11:8]<=7;data[445][7:5]<=4;data[445][4:0]<=1;
			data[446][11:8]<=9;data[446][7:5]<=4;data[446][4:0]<=1;
			data[447][11:8]<=11;data[447][7:5]<=4;data[447][4:0]<=1;
			data[448][11:8]<=7;data[448][7:5]<=4;data[448][4:0]<=2;
			data[449][11:8]<=11;data[449][7:5]<=4;data[449][4:0]<=1;
			data[450][11:8]<=9;data[450][7:5]<=4;data[450][4:0]<=1;
			data[451][11:8]<=11;data[451][7:5]<=4;data[451][4:0]<=2;
			data[452][11:8]<=13;data[452][7:5]<=4;data[452][4:0]<=1;
			data[453][11:8]<=2;data[453][7:5]<=3;data[453][4:0]<=1;
			data[454][11:8]<=9;data[454][7:5]<=4;data[454][4:0]<=1;
			data[455][11:8]<=11;data[455][7:5]<=4;data[455][4:0]<=1;
			data[456][11:8]<=13;data[456][7:5]<=4;data[456][4:0]<=1;
			data[457][11:8]<=2;data[457][7:5]<=3;data[457][4:0]<=1;
			data[458][11:8]<=4;data[458][7:5]<=3;data[458][4:0]<=1;
			data[459][11:8]<=6;data[459][7:5]<=3;data[459][4:0]<=1;
			data[460][11:8]<=7;data[460][7:5]<=3;data[460][4:0]<=1;
			data[461][11:8]<=9;data[461][7:5]<=3;data[461][4:0]<=1;
			data[462][11:8]<=6;data[462][7:5]<=3;data[462][4:0]<=2;
			data[463][11:8]<=2;data[463][7:5]<=3;data[463][4:0]<=1;
			data[464][11:8]<=4;data[464][7:5]<=3;data[464][4:0]<=1;
			data[465][11:8]<=6;data[465][7:5]<=3;data[465][4:0]<=2;
			data[466][11:8]<=4;data[466][7:5]<=3;data[466][4:0]<=1;
			data[467][11:8]<=2;data[467][7:5]<=3;data[467][4:0]<=1;
			data[468][11:8]<=4;data[468][7:5]<=3;data[468][4:0]<=1;
			data[469][11:8]<=13;data[469][7:5]<=4;data[469][4:0]<=1;
			data[470][11:8]<=2;data[470][7:5]<=3;data[470][4:0]<=1;
			data[471][11:8]<=4;data[471][7:5]<=3;data[471][4:0]<=1;
			data[472][11:8]<=6;data[472][7:5]<=3;data[472][4:0]<=1;
			data[473][11:8]<=4;data[473][7:5]<=3;data[473][4:0]<=1;
			data[474][11:8]<=2;data[474][7:5]<=3;data[474][4:0]<=1;
			data[475][11:8]<=13;data[475][7:5]<=4;data[475][4:0]<=1;
			data[476][11:8]<=2;data[476][7:5]<=3;data[476][4:0]<=2;
			data[477][11:8]<=11;data[477][7:5]<=4;data[477][4:0]<=1;
			data[478][11:8]<=13;data[478][7:5]<=4;data[478][4:0]<=1;
			data[479][11:8]<=2;data[479][7:5]<=3;data[479][4:0]<=2;
			data[480][11:8]<=2;data[480][7:5]<=4;data[480][4:0]<=1;
			data[481][11:8]<=4;data[481][7:5]<=4;data[481][4:0]<=1;
			data[482][11:8]<=6;data[482][7:5]<=4;data[482][4:0]<=1;
			data[483][11:8]<=7;data[483][7:5]<=4;data[483][4:0]<=1;
			data[484][11:8]<=6;data[484][7:5]<=4;data[484][4:0]<=1;
			data[485][11:8]<=4;data[485][7:5]<=4;data[485][4:0]<=1;
			data[486][11:8]<=6;data[486][7:5]<=4;data[486][4:0]<=1;
			data[487][11:8]<=2;data[487][7:5]<=3;data[487][4:0]<=1;
			data[488][11:8]<=13;data[488][7:5]<=4;data[488][4:0]<=1;
			data[489][11:8]<=2;data[489][7:5]<=3;data[489][4:0]<=1;
			data[490][11:8]<=11;data[490][7:5]<=4;data[490][4:0]<=2;
			data[491][11:8]<=2;data[491][7:5]<=3;data[491][4:0]<=1;
			data[492][11:8]<=13;data[492][7:5]<=4;data[492][4:0]<=1;
			data[493][11:8]<=11;data[493][7:5]<=4;data[493][4:0]<=2;
			data[494][11:8]<=9;data[494][7:5]<=4;data[494][4:0]<=1;
			data[495][11:8]<=7;data[495][7:5]<=4;data[495][4:0]<=1;
			data[496][11:8]<=9;data[496][7:5]<=4;data[496][4:0]<=1;
			data[497][11:8]<=7;data[497][7:5]<=4;data[497][4:0]<=1;
			data[498][11:8]<=6;data[498][7:5]<=4;data[498][4:0]<=1;
			data[499][11:8]<=7;data[499][7:5]<=4;data[499][4:0]<=1;
			data[500][11:8]<=9;data[500][7:5]<=4;data[500][4:0]<=1;
			data[501][11:8]<=11;data[501][7:5]<=4;data[501][4:0]<=1;
			data[502][11:8]<=13;data[502][7:5]<=4;data[502][4:0]<=1;
			data[503][11:8]<=2;data[503][7:5]<=4;data[503][4:0]<=1;
			data[504][11:8]<=11;data[504][7:5]<=4;data[504][4:0]<=2;
			data[505][11:8]<=2;data[505][7:5]<=3;data[505][4:0]<=1;
			data[506][11:8]<=13;data[506][7:5]<=4;data[506][4:0]<=1;
			data[507][11:8]<=2;data[507][7:5]<=3;data[507][4:0]<=2;
			data[508][11:8]<=13;data[508][7:5]<=4;data[508][4:0]<=1;
			data[509][11:8]<=11;data[509][7:5]<=4;data[509][4:0]<=1;
			data[510][11:8]<=13;data[510][7:5]<=4;data[510][4:0]<=1;
			data[511][11:8]<=2;data[511][7:5]<=3;data[511][4:0]<=1;
			data[512][11:8]<=4;data[512][7:5]<=3;data[512][4:0]<=1;
			data[513][11:8]<=2;data[513][7:5]<=3;data[513][4:0]<=1;
			data[514][11:8]<=13;data[514][7:5]<=4;data[514][4:0]<=1;
			data[515][11:8]<=2;data[515][7:5]<=3;data[515][4:0]<=1;
			data[516][11:8]<=11;data[516][7:5]<=4;data[516][4:0]<=1;
			data[517][11:8]<=13;data[517][7:5]<=4;data[517][4:0]<=1;
			data[518][11:8]<=6;data[518][7:5]<=3;data[518][4:0]<=2;
			data[519][11:8]<=6;data[519][7:5]<=4;data[519][4:0]<=2;
			data[520][11:8]<=7;data[520][7:5]<=4;data[520][4:0]<=2;
			data[521][11:8]<=6;data[521][7:5]<=4;data[521][4:0]<=2;
			data[522][11:8]<=4;data[522][7:5]<=4;data[522][4:0]<=2;
			data[523][11:8]<=4;data[523][7:5]<=3;data[523][4:0]<=2;
			data[524][11:8]<=6;data[524][7:5]<=3;data[524][4:0]<=2;
			data[525][11:8]<=4;data[525][7:5]<=3;data[525][4:0]<=2;
			data[526][11:8]<=2;data[526][7:5]<=3;data[526][4:0]<=2;
			data[527][11:8]<=6;data[527][7:5]<=4;data[527][4:0]<=2;
			data[528][11:8]<=2;data[528][7:5]<=4;data[528][4:0]<=2;
			data[529][11:8]<=11;data[529][7:5]<=4;data[529][4:0]<=2;
			data[530][11:8]<=9;data[530][7:5]<=4;data[530][4:0]<=2;
			data[531][11:8]<=9;data[531][7:5]<=5;data[531][4:0]<=2;
			data[532][11:8]<=7;data[532][7:5]<=5;data[532][4:0]<=2;
			data[533][11:8]<=9;data[533][7:5]<=5;data[533][4:0]<=2;
			data[534][11:8]<=11;data[534][7:5]<=5;data[534][4:0]<=2;
			data[535][11:8]<=11;data[535][7:5]<=4;data[535][4:0]<=2;
			data[536][11:8]<=13;data[536][7:5]<=4;data[536][4:0]<=2;
			data[537][11:8]<=11;data[537][7:5]<=4;data[537][4:0]<=2;
			data[538][11:8]<=13;data[538][7:5]<=4;data[538][4:0]<=2;
			data[539][11:8]<=9;data[539][7:5]<=5;data[539][4:0]<=2;
			data[540][11:8]<=7;data[540][7:5]<=5;data[540][4:0]<=2;
			data[541][11:8]<=9;data[541][7:5]<=5;data[541][4:0]<=2;
			data[542][11:8]<=11;data[542][7:5]<=5;data[542][4:0]<=2;
			data[543][11:8]<=11;data[543][7:5]<=4;data[543][4:0]<=2;
			data[544][11:8]<=9;data[544][7:5]<=4;data[544][4:0]<=2;
			data[545][11:8]<=11;data[545][7:5]<=4;data[545][4:0]<=2;
			data[546][11:8]<=13;data[546][7:5]<=4;data[546][4:0]<=2;
			data[547][11:8]<=13;data[547][7:5]<=4;data[547][4:0]<=2;
			data[548][11:8]<=11;data[548][7:5]<=4;data[548][4:0]<=2;
			data[549][11:8]<=13;data[549][7:5]<=4;data[549][4:0]<=2;
			data[550][11:8]<=2;data[550][7:5]<=4;data[550][4:0]<=2;
			data[551][11:8]<=2;data[551][7:5]<=3;data[551][4:0]<=2;
			data[552][11:8]<=4;data[552][7:5]<=3;data[552][4:0]<=2;
			data[553][11:8]<=2;data[553][7:5]<=3;data[553][4:0]<=2;
			data[554][11:8]<=13;data[554][7:5]<=4;data[554][4:0]<=2;
			data[555][11:8]<=13;data[555][7:5]<=5;data[555][4:0]<=2;
			data[556][11:8]<=2;data[556][7:5]<=4;data[556][4:0]<=2;
			data[557][11:8]<=13;data[557][7:5]<=5;data[557][4:0]<=2;
			data[558][11:8]<=11;data[558][7:5]<=5;data[558][4:0]<=2;
			data[559][11:8]<=11;data[559][7:5]<=4;data[559][4:0]<=2;
			data[560][11:8]<=9;data[560][7:5]<=4;data[560][4:0]<=2;
			data[561][11:8]<=11;data[561][7:5]<=4;data[561][4:0]<=2;
			data[562][11:8]<=13;data[562][7:5]<=4;data[562][4:0]<=2;
			data[563][11:8]<=13;data[563][7:5]<=5;data[563][4:0]<=2;
			data[564][11:8]<=6;data[564][7:5]<=4;data[564][4:0]<=2;
			data[565][11:8]<=4;data[565][7:5]<=4;data[565][4:0]<=2;
			data[566][11:8]<=2;data[566][7:5]<=4;data[566][4:0]<=2;
			data[567][11:8]<=2;data[567][7:5]<=3;data[567][4:0]<=2;
			data[568][11:8]<=4;data[568][7:5]<=3;data[568][4:0]<=2;
			data[569][11:8]<=7;data[569][7:5]<=3;data[569][4:0]<=2;
			data[570][11:8]<=6;data[570][7:5]<=3;data[570][4:0]<=2;
			data[571][11:8]<=6;data[571][7:5]<=4;data[571][4:0]<=2;
			data[572][11:8]<=9;data[572][7:5]<=4;data[572][4:0]<=2;
			data[573][11:8]<=6;data[573][7:5]<=3;data[573][4:0]<=2;
			data[574][11:8]<=2;data[574][7:5]<=3;data[574][4:0]<=2;
			data[575][11:8]<=7;data[575][7:5]<=3;data[575][4:0]<=2;
			data[576][11:8]<=6;data[576][7:5]<=3;data[576][4:0]<=2;
			data[577][11:8]<=7;data[577][7:5]<=3;data[577][4:0]<=2;
			data[578][11:8]<=4;data[578][7:5]<=3;data[578][4:0]<=2;
			data[579][11:8]<=9;data[579][7:5]<=4;data[579][4:0]<=2;
			data[580][11:8]<=7;data[580][7:5]<=4;data[580][4:0]<=2;
			data[581][11:8]<=9;data[581][7:5]<=4;data[581][4:0]<=2;
			data[582][11:8]<=6;data[582][7:5]<=4;data[582][4:0]<=2;
			data[583][11:8]<=2;data[583][7:5]<=3;data[583][4:0]<=1;
			data[584][11:8]<=13;data[584][7:5]<=4;data[584][4:0]<=1;
			data[585][11:8]<=2;data[585][7:5]<=3;data[585][4:0]<=2;
			data[586][11:8]<=6;data[586][7:5]<=4;data[586][4:0]<=2;
			data[587][11:8]<=9;data[587][7:5]<=4;data[587][4:0]<=2;
			data[588][11:8]<=9;data[588][7:5]<=4;data[588][4:0]<=1;
			data[589][11:8]<=11;data[589][7:5]<=4;data[589][4:0]<=1;
			data[590][11:8]<=13;data[590][7:5]<=4;data[590][4:0]<=2;
			data[591][11:8]<=9;data[591][7:5]<=4;data[591][4:0]<=2;
			data[592][11:8]<=6;data[592][7:5]<=4;data[592][4:0]<=2;
			data[593][11:8]<=2;data[593][7:5]<=3;data[593][4:0]<=1;
			data[594][11:8]<=4;data[594][7:5]<=3;data[594][4:0]<=1;
			data[595][11:8]<=6;data[595][7:5]<=3;data[595][4:0]<=2;
			data[596][11:8]<=2;data[596][7:5]<=3;data[596][4:0]<=2;
			data[597][11:8]<=6;data[597][7:5]<=3;data[597][4:0]<=2;
			data[598][11:8]<=6;data[598][7:5]<=3;data[598][4:0]<=1;
			data[599][11:8]<=4;data[599][7:5]<=3;data[599][4:0]<=1;
			data[600][11:8]<=2;data[600][7:5]<=3;data[600][4:0]<=2;
			data[601][11:8]<=13;data[601][7:5]<=4;data[601][4:0]<=2;
			data[602][11:8]<=11;data[602][7:5]<=4;data[602][4:0]<=2;
			data[603][11:8]<=11;data[603][7:5]<=4;data[603][4:0]<=1;
			data[604][11:8]<=9;data[604][7:5]<=4;data[604][4:0]<=1;
			data[605][11:8]<=11;data[605][7:5]<=4;data[605][4:0]<=2;
			data[606][11:8]<=13;data[606][7:5]<=4;data[606][4:0]<=2;
			data[607][11:8]<=2;data[607][7:5]<=3;data[607][4:0]<=2;
			data[608][11:8]<=6;data[608][7:5]<=3;data[608][4:0]<=1;
			data[609][11:8]<=4;data[609][7:5]<=3;data[609][4:0]<=1;
			data[610][11:8]<=2;data[610][7:5]<=3;data[610][4:0]<=2;
			data[611][11:8]<=6;data[611][7:5]<=3;data[611][4:0]<=2;
			data[612][11:8]<=7;data[612][7:5]<=4;data[612][4:0]<=2;
			data[613][11:8]<=2;data[613][7:5]<=4;data[613][4:0]<=1;
			data[614][11:8]<=13;data[614][7:5]<=4;data[614][4:0]<=1;
			data[615][11:8]<=11;data[615][7:5]<=4;data[615][4:0]<=2;
			data[616][11:8]<=11;data[616][7:5]<=4;data[616][4:0]<=2;
			data[617][11:8]<=9;data[617][7:5]<=4;data[617][4:0]<=2;
			data[618][11:8]<=4;data[618][7:5]<=4;data[618][4:0]<=2;
			data[619][11:8]<=9;data[619][7:5]<=4;data[619][4:0]<=2;
			data[620][11:8]<=9;data[620][7:5]<=4;data[620][4:0]<=2;
			data[621][11:8]<=6;data[621][7:5]<=4;data[621][4:0]<=6;
			data[622][11:8]<=6;data[622][7:5]<=3;data[622][4:0]<=2;
			data[623][11:8]<=6;data[623][7:5]<=3;data[623][4:0]<=2;
			data[624][11:8]<=7;data[624][7:5]<=3;data[624][4:0]<=2;
			data[625][11:8]<=6;data[625][7:5]<=3;data[625][4:0]<=2;
			data[626][11:8]<=4;data[626][7:5]<=3;data[626][4:0]<=2;
			data[627][11:8]<=2;data[627][7:5]<=3;data[627][4:0]<=6;
			data[628][11:8]<=2;data[628][7:5]<=3;data[628][4:0]<=2;
			data[629][11:8]<=2;data[629][7:5]<=3;data[629][4:0]<=2;
			data[630][11:8]<=4;data[630][7:5]<=3;data[630][4:0]<=2;
			data[631][11:8]<=2;data[631][7:5]<=3;data[631][4:0]<=2;
			data[632][11:8]<=13;data[632][7:5]<=4;data[632][4:0]<=2;
			data[633][11:8]<=11;data[633][7:5]<=4;data[633][4:0]<=8;
			data[634][11:8]<=2;data[634][7:5]<=3;data[634][4:0]<=8;
			data[635][11:8]<=2;data[635][7:5]<=3;data[635][4:0]<=2;
			data[636][11:8]<=12;data[636][7:5]<=4;data[636][4:0]<=2;
			data[637][11:8]<=11;data[637][7:5]<=4;data[637][4:0]<=2;
			data[638][11:8]<=12;data[638][7:5]<=4;data[638][4:0]<=2;
			data[639][11:8]<=9;data[639][7:5]<=4;data[639][4:0]<=6;
			data[640][11:8]<=9;data[640][7:5]<=4;data[640][4:0]<=2;
			data[641][11:8]<=9;data[641][7:5]<=4;data[641][4:0]<=6;
			data[642][11:8]<=9;data[642][7:5]<=4;data[642][4:0]<=2;
			data[643][11:8]<=9;data[643][7:5]<=4;data[643][4:0]<=2;
			data[644][11:8]<=11;data[644][7:5]<=4;data[644][4:0]<=2;
			data[645][11:8]<=9;data[645][7:5]<=4;data[645][4:0]<=2;
			data[646][11:8]<=7;data[646][7:5]<=4;data[646][4:0]<=2;
			data[647][11:8]<=6;data[647][7:5]<=4;data[647][4:0]<=6;
			data[648][11:8]<=6;data[648][7:5]<=4;data[648][4:0]<=2;
			data[649][11:8]<=6;data[649][7:5]<=4;data[649][4:0]<=2;
			data[650][11:8]<=7;data[650][7:5]<=4;data[650][4:0]<=2;
			data[651][11:8]<=6;data[651][7:5]<=4;data[651][4:0]<=2;
			data[652][11:8]<=4;data[652][7:5]<=4;data[652][4:0]<=2;
			data[653][11:8]<=2;data[653][7:5]<=3;data[653][4:0]<=2;
			data[654][11:8]<=12;data[654][7:5]<=4;data[654][4:0]<=2;
			data[655][11:8]<=11;data[655][7:5]<=4;data[655][4:0]<=2;
			data[656][11:8]<=12;data[656][7:5]<=4;data[656][4:0]<=2;
			data[657][11:8]<=9;data[657][7:5]<=4;data[657][4:0]<=6;
			data[658][11:8]<=9;data[658][7:5]<=4;data[658][4:0]<=2;
			data[659][11:8]<=7;data[659][7:5]<=4;data[659][4:0]<=4;
			data[660][11:8]<=2;data[660][7:5]<=3;data[660][4:0]<=4;
			data[661][11:8]<=13;data[661][7:5]<=4;data[661][4:0]<=6;
			data[662][11:8]<=13;data[662][7:5]<=4;data[662][4:0]<=2;
			data[663][11:8]<=9;data[663][7:5]<=3;data[663][4:0]<=8;
			data[664][11:8]<=9;data[664][7:5]<=4;data[664][4:0]<=6;
			data[665][11:8]<=7;data[665][7:5]<=4;data[665][4:0]<=2;
			data[666][11:8]<=6;data[666][7:5]<=3;data[666][4:0]<=8;
			data[667][11:8]<=6;data[667][7:5]<=3;data[667][4:0]<=6;
			data[668][11:8]<=4;data[668][7:5]<=3;data[668][4:0]<=2;
			data[669][11:8]<=2;data[669][7:5]<=3;data[669][4:0]<=12;
			data[670][11:8]<=2;data[670][7:5]<=4;data[670][4:0]<=4;
			data[671][11:8]<=2;data[671][7:5]<=3;data[671][4:0]<=8;
			data[672][11:8]<=13;data[672][7:5]<=4;data[672][4:0]<=8;
			data[673][11:8]<=2;data[673][7:5]<=3;data[673][4:0]<=4;
			data[674][11:8]<=2;data[674][7:5]<=4;data[674][4:0]<=4;
			data[675][11:8]<=13;data[675][7:5]<=5;data[675][4:0]<=4;
			data[676][11:8]<=13;data[676][7:5]<=4;data[676][4:0]<=4;
			data[677][11:8]<=11;data[677][7:5]<=4;data[677][4:0]<=4;
			data[678][11:8]<=11;data[678][7:5]<=5;data[678][4:0]<=4;
			data[679][11:8]<=9;data[679][7:5]<=5;data[679][4:0]<=4;
			data[680][11:8]<=9;data[680][7:5]<=4;data[680][4:0]<=4;
			data[681][11:8]<=7;data[681][7:5]<=4;data[681][4:0]<=4;
			data[682][11:8]<=7;data[682][7:5]<=3;data[682][4:0]<=4;
			data[683][11:8]<=6;data[683][7:5]<=3;data[683][4:0]<=4;
			data[684][11:8]<=6;data[684][7:5]<=4;data[684][4:0]<=4;
			data[685][11:8]<=4;data[685][7:5]<=4;data[685][4:0]<=4;
			data[686][11:8]<=11;data[686][7:5]<=4;data[686][4:0]<=4;
			data[687][11:8]<=4;data[687][7:5]<=4;data[687][4:0]<=4;
			data[688][11:8]<=4;data[688][7:5]<=3;data[688][4:0]<=4;
			data[689][11:8]<=6;data[689][7:5]<=3;data[689][4:0]<=4;
			data[690][11:8]<=6;data[690][7:5]<=4;data[690][4:0]<=4;
			data[691][11:8]<=4;data[691][7:5]<=4;data[691][4:0]<=4;
			data[692][11:8]<=4;data[692][7:5]<=3;data[692][4:0]<=4;
			data[693][11:8]<=2;data[693][7:5]<=3;data[693][4:0]<=4;
			data[694][11:8]<=2;data[694][7:5]<=4;data[694][4:0]<=4;
			data[695][11:8]<=13;data[695][7:5]<=5;data[695][4:0]<=4;
			data[696][11:8]<=13;data[696][7:5]<=4;data[696][4:0]<=4;
			data[697][11:8]<=11;data[697][7:5]<=4;data[697][4:0]<=4;
			data[698][11:8]<=11;data[698][7:5]<=3;data[698][4:0]<=4;
			data[699][11:8]<=9;data[699][7:5]<=3;data[699][4:0]<=4;
			data[700][11:8]<=9;data[700][7:5]<=4;data[700][4:0]<=4;
			data[701][11:8]<=7;data[701][7:5]<=4;data[701][4:0]<=6;
			data[702][11:8]<=4;data[702][7:5]<=3;data[702][4:0]<=2;
			data[703][11:8]<=9;data[703][7:5]<=4;data[703][4:0]<=4;
			data[704][11:8]<=4;data[704][7:5]<=3;data[704][4:0]<=4;
			data[705][11:8]<=6;data[705][7:5]<=3;data[705][4:0]<=8;
			data[706][11:8]<=0;data[706][7:5]<=4;data[706][4:0]<=4;
			data[707][11:8]<=0;data[707][7:5]<=4;data[707][4:0]<=4;

			data[711][11:8]<=11;data[711][7:5]<=4;data[711][4:0]<=8;
			data[712][11:8]<=2;data[712][7:5]<=3;data[712][4:0]<=4;
			data[713][11:8]<=4;data[713][7:5]<=3;data[713][4:0]<=4;
			data[714][11:8]<=11;data[714][7:5]<=4;data[714][4:0]<=8;
			data[715][11:8]<=2;data[715][7:5]<=3;data[715][4:0]<=4;
			data[716][11:8]<=4;data[716][7:5]<=3;data[716][4:0]<=4;
			data[717][11:8]<=6;data[717][7:5]<=3;data[717][4:0]<=8;
			data[718][11:8]<=9;data[718][7:5]<=3;data[718][4:0]<=4;
			data[719][11:8]<=11;data[719][7:5]<=3;data[719][4:0]<=4;
			data[720][11:8]<=4;data[720][7:5]<=3;data[720][4:0]<=8;
			data[721][11:8]<=2;data[721][7:5]<=3;data[721][4:0]<=4;
			data[722][11:8]<=13;data[722][7:5]<=4;data[722][4:0]<=4;
			data[723][11:8]<=11;data[723][7:5]<=4;data[723][4:0]<=12;
			data[724][11:8]<=9;data[724][7:5]<=4;data[724][4:0]<=4;
			data[725][11:8]<=2;data[725][7:5]<=3;data[725][4:0]<=8;
			data[726][11:8]<=13;data[726][7:5]<=4;data[726][4:0]<=6;
			data[727][11:8]<=4;data[727][7:5]<=3;data[727][4:0]<=2;
			data[728][11:8]<=11;data[728][7:5]<=4;data[728][4:0]<=16;
			data[729][11:8]<=0;data[729][7:5]<=4;data[729][4:0]<=16;
			data[730][11:8]<=0;data[730][7:5]<=4;data[730][4:0]<=2;
			data[731][11:8]<=11;data[731][7:5]<=4;data[731][4:0]<=2;
			data[732][11:8]<=6;data[732][7:5]<=3;data[732][4:0]<=2;
			data[733][11:8]<=4;data[733][7:5]<=3;data[733][4:0]<=2;
			data[734][11:8]<=6;data[734][7:5]<=3;data[734][4:0]<=4;
			data[735][11:8]<=2;data[735][7:5]<=3;data[735][4:0]<=4;
			data[736][11:8]<=13;data[736][7:5]<=4;data[736][4:0]<=4;
			data[737][11:8]<=2;data[737][7:5]<=3;data[737][4:0]<=2;
			data[738][11:8]<=4;data[738][7:5]<=3;data[738][4:0]<=4;
			data[739][11:8]<=13;data[739][7:5]<=4;data[739][4:0]<=6;
			data[740][11:8]<=0;data[740][7:5]<=4;data[740][4:0]<=2;
			data[741][11:8]<=11;data[741][7:5]<=4;data[741][4:0]<=2;
			data[742][11:8]<=6;data[742][7:5]<=3;data[742][4:0]<=2;
			data[743][11:8]<=4;data[743][7:5]<=3;data[743][4:0]<=2;
			data[744][11:8]<=6;data[744][7:5]<=3;data[744][4:0]<=4;
			data[745][11:8]<=2;data[745][7:5]<=3;data[745][4:0]<=4;
			data[746][11:8]<=13;data[746][7:5]<=4;data[746][4:0]<=4;
			data[747][11:8]<=2;data[747][7:5]<=3;data[747][4:0]<=2;
			data[748][11:8]<=4;data[748][7:5]<=3;data[748][4:0]<=4;
			data[749][11:8]<=13;data[749][7:5]<=4;data[749][4:0]<=4;
			data[750][11:8]<=11;data[750][7:5]<=4;data[750][4:0]<=12;
			data[751][11:8]<=9;data[751][7:5]<=4;data[751][4:0]<=2;
			data[752][11:8]<=2;data[752][7:5]<=3;data[752][4:0]<=2;
			data[753][11:8]<=13;data[753][7:5]<=4;data[753][4:0]<=10;
			data[754][11:8]<=13;data[754][7:5]<=4;data[754][4:0]<=2;
			data[755][11:8]<=2;data[755][7:5]<=3;data[755][4:0]<=2;
			data[756][11:8]<=4;data[756][7:5]<=3;data[756][4:0]<=2;
			data[757][11:8]<=11;data[757][7:5]<=4;data[757][4:0]<=4;
			data[758][11:8]<=11;data[758][7:5]<=4;data[758][4:0]<=14;
			data[759][11:8]<=2;data[759][7:5]<=3;data[759][4:0]<=4;
			data[760][11:8]<=2;data[760][7:5]<=2;data[760][4:0]<=4;
			data[761][11:8]<=13;data[761][7:5]<=3;data[761][4:0]<=4;
			data[762][11:8]<=2;data[762][7:5]<=2;data[762][4:0]<=4;
			data[763][11:8]<=9;data[763][7:5]<=3;data[763][4:0]<=3;
			data[764][11:8]<=2;data[764][7:5]<=3;data[764][4:0]<=3;
			data[765][11:8]<=11;data[765][7:5]<=3;data[765][4:0]<=4;
			data[766][11:8]<=9;data[766][7:5]<=3;data[766][4:0]<=8;
			data[767][11:8]<=2;data[767][7:5]<=3;data[767][4:0]<=2;
			data[768][11:8]<=2;data[768][7:5]<=2;data[768][4:0]<=2;
			data[769][11:8]<=13;data[769][7:5]<=3;data[769][4:0]<=4;
			data[770][11:8]<=2;data[770][7:5]<=2;data[770][4:0]<=4;
			data[771][11:8]<=9;data[771][7:5]<=3;data[771][4:0]<=3;
			data[772][11:8]<=6;data[772][7:5]<=3;data[772][4:0]<=3;
			data[773][11:8]<=11;data[773][7:5]<=3;data[773][4:0]<=2;
			data[774][11:8]<=11;data[774][7:5]<=3;data[774][4:0]<=2;
			data[775][11:8]<=13;data[775][7:5]<=3;data[775][4:0]<=2;
			data[776][11:8]<=9;data[776][7:5]<=3;data[776][4:0]<=8;
			data[777][11:8]<=9;data[777][7:5]<=3;data[777][4:0]<=2;
			data[778][11:8]<=9;data[778][7:5]<=3;data[778][4:0]<=2;
			data[779][11:8]<=7;data[779][7:5]<=3;data[779][4:0]<=2;
			data[780][11:8]<=7;data[780][7:5]<=3;data[780][4:0]<=2;
			data[781][11:8]<=6;data[781][7:5]<=3;data[781][4:0]<=2;
			data[782][11:8]<=6;data[782][7:5]<=3;data[782][4:0]<=3;
			data[783][11:8]<=2;data[783][7:5]<=3;data[783][4:0]<=3;
			data[784][11:8]<=11;data[784][7:5]<=4;data[784][4:0]<=2;
			data[785][11:8]<=4;data[785][7:5]<=3;data[785][4:0]<=2;
			data[786][11:8]<=2;data[786][7:5]<=3;data[786][4:0]<=6;
			data[787][11:8]<=2;data[787][7:5]<=3;data[787][4:0]<=4;
			data[788][11:8]<=9;data[788][7:5]<=3;data[788][4:0]<=2;
			data[789][11:8]<=9;data[789][7:5]<=3;data[789][4:0]<=2;
			data[790][11:8]<=7;data[790][7:5]<=3;data[790][4:0]<=2;
			data[791][11:8]<=7;data[791][7:5]<=3;data[791][4:0]<=2;
			data[792][11:8]<=6;data[792][7:5]<=3;data[792][4:0]<=2;
			data[793][11:8]<=6;data[793][7:5]<=3;data[793][4:0]<=3;
			data[794][11:8]<=4;data[794][7:5]<=3;data[794][4:0]<=3;
			data[795][11:8]<=2;data[795][7:5]<=3;data[795][4:0]<=4;
			data[796][11:8]<=4;data[796][7:5]<=3;data[796][4:0]<=10;
			data[797][11:8]<=2;data[797][7:5]<=3;data[797][4:0]<=4;
			data[798][11:8]<=2;data[798][7:5]<=2;data[798][4:0]<=2;
			data[799][11:8]<=13;data[799][7:5]<=3;data[799][4:0]<=4;
			data[800][11:8]<=2;data[800][7:5]<=2;data[800][4:0]<=4;
			data[801][11:8]<=9;data[801][7:5]<=3;data[801][4:0]<=3;
			data[802][11:8]<=6;data[802][7:5]<=3;data[802][4:0]<=3;
			data[803][11:8]<=11;data[803][7:5]<=3;data[803][4:0]<=4;
			data[804][11:8]<=9;data[804][7:5]<=3;data[804][4:0]<=10;
			data[805][11:8]<=2;data[805][7:5]<=3;data[805][4:0]<=2;
			data[806][11:8]<=2;data[806][7:5]<=2;data[806][4:0]<=2;
			data[807][11:8]<=13;data[807][7:5]<=3;data[807][4:0]<=4;
			data[808][11:8]<=2;data[808][7:5]<=2;data[808][4:0]<=4;
			data[809][11:8]<=4;data[809][7:5]<=2;data[809][4:0]<=3;
			data[810][11:8]<=9;data[810][7:5]<=3;data[810][4:0]<=3;
			data[811][11:8]<=4;data[811][7:5]<=2;data[811][4:0]<=2;
			data[812][11:8]<=4;data[812][7:5]<=2;data[812][4:0]<=3;
			data[813][11:8]<=6;data[813][7:5]<=2;data[813][4:0]<=10;
			data[814][11:8]<=9;data[814][7:5]<=3;data[814][4:0]<=10;
			data[815][11:8]<=7;data[815][7:5]<=3;data[815][4:0]<=2;
			data[816][11:8]<=6;data[816][7:5]<=3;data[816][4:0]<=2;
			data[817][11:8]<=7;data[817][7:5]<=3;data[817][4:0]<=2;
			data[818][11:8]<=9;data[818][7:5]<=3;data[818][4:0]<=3;
			data[819][11:8]<=2;data[819][7:5]<=3;data[819][4:0]<=2;
			data[820][11:8]<=9;data[820][7:5]<=3;data[820][4:0]<=3;
			data[821][11:8]<=11;data[821][7:5]<=3;data[821][4:0]<=3;
			data[822][11:8]<=13;data[822][7:5]<=3;data[822][4:0]<=2;
			data[823][11:8]<=2;data[823][7:5]<=2;data[823][4:0]<=2;
			data[824][11:8]<=13;data[824][7:5]<=3;data[824][4:0]<=2;
			data[825][11:8]<=9;data[825][7:5]<=3;data[825][4:0]<=3;
			data[826][11:8]<=6;data[826][7:5]<=3;data[826][4:0]<=4;
			data[827][11:8]<=6;data[827][7:5]<=3;data[827][4:0]<=4;
			data[828][11:8]<=4;data[828][7:5]<=3;data[828][4:0]<=2;
			data[829][11:8]<=4;data[829][7:5]<=3;data[829][4:0]<=12;
			data[830][11:8]<=9;data[830][7:5]<=4;data[830][4:0]<=4;
			data[831][11:8]<=11;data[831][7:5]<=4;data[831][4:0]<=4;
			data[832][11:8]<=2;data[832][7:5]<=3;data[832][4:0]<=4;
			data[833][11:8]<=4;data[833][7:5]<=3;data[833][4:0]<=2;
			data[834][11:8]<=9;data[834][7:5]<=4;data[834][4:0]<=2;
			data[835][11:8]<=9;data[835][7:5]<=4;data[835][4:0]<=4;
			data[836][11:8]<=11;data[836][7:5]<=4;data[836][4:0]<=4;
			data[837][11:8]<=2;data[837][7:5]<=3;data[837][4:0]<=2;
			data[838][11:8]<=4;data[838][7:5]<=3;data[838][4:0]<=2;
			data[839][11:8]<=9;data[839][7:5]<=4;data[839][4:0]<=4;
			data[840][11:8]<=6;data[840][7:5]<=3;data[840][4:0]<=4;
			data[841][11:8]<=4;data[841][7:5]<=3;data[841][4:0]<=4;
			data[842][11:8]<=4;data[842][7:5]<=3;data[842][4:0]<=4;
			data[843][11:8]<=2;data[843][7:5]<=3;data[843][4:0]<=2;
			data[844][11:8]<=13;data[844][7:5]<=4;data[844][4:0]<=2;
			data[845][11:8]<=13;data[845][7:5]<=4;data[845][4:0]<=4;
			data[846][11:8]<=2;data[846][7:5]<=3;data[846][4:0]<=4;
			data[847][11:8]<=13;data[847][7:5]<=4;data[847][4:0]<=4;
			data[848][11:8]<=9;data[848][7:5]<=4;data[848][4:0]<=4;
			data[849][11:8]<=9;data[849][7:5]<=4;data[849][4:0]<=4;
			data[850][11:8]<=11;data[850][7:5]<=4;data[850][4:0]<=4;
			data[851][11:8]<=2;data[851][7:5]<=3;data[851][4:0]<=4;
			data[852][11:8]<=4;data[852][7:5]<=3;data[852][4:0]<=2;
			data[853][11:8]<=9;data[853][7:5]<=4;data[853][4:0]<=2;
			data[854][11:8]<=9;data[854][7:5]<=4;data[854][4:0]<=4;
			data[855][11:8]<=11;data[855][7:5]<=4;data[855][4:0]<=4;
			data[856][11:8]<=2;data[856][7:5]<=3;data[856][4:0]<=2;
			data[857][11:8]<=4;data[857][7:5]<=3;data[857][4:0]<=2;
			data[858][11:8]<=9;data[858][7:5]<=4;data[858][4:0]<=4;
			data[859][11:8]<=6;data[859][7:5]<=3;data[859][4:0]<=4;
			data[860][11:8]<=4;data[860][7:5]<=3;data[860][4:0]<=4;
			data[861][11:8]<=4;data[861][7:5]<=3;data[861][4:0]<=4;
			data[862][11:8]<=2;data[862][7:5]<=3;data[862][4:0]<=2;
			data[863][11:8]<=13;data[863][7:5]<=4;data[863][4:0]<=2;
			data[864][11:8]<=13;data[864][7:5]<=4;data[864][4:0]<=4;
			data[865][11:8]<=2;data[865][7:5]<=3;data[865][4:0]<=8;
			data[866][11:8]<=9;data[866][7:5]<=3;data[866][4:0]<=2;
			data[867][11:8]<=11;data[867][7:5]<=3;data[867][4:0]<=2;
			data[868][11:8]<=9;data[868][7:5]<=3;data[868][4:0]<=3;
			data[869][11:8]<=6;data[869][7:5]<=3;data[869][4:0]<=2;
			data[870][11:8]<=9;data[870][7:5]<=3;data[870][4:0]<=3;
			data[871][11:8]<=2;data[871][7:5]<=3;data[871][4:0]<=2;
			data[872][11:8]<=2;data[872][7:5]<=3;data[872][4:0]<=2;
			data[873][11:8]<=4;data[873][7:5]<=3;data[873][4:0]<=2;
			data[874][11:8]<=6;data[874][7:5]<=3;data[874][4:0]<=2;
			data[875][11:8]<=11;data[875][7:5]<=3;data[875][4:0]<=2;
			data[876][11:8]<=9;data[876][7:5]<=3;data[876][4:0]<=4;
			data[877][11:8]<=6;data[877][7:5]<=3;data[877][4:0]<=2;
			data[878][11:8]<=9;data[878][7:5]<=3;data[878][4:0]<=2;
			data[879][11:8]<=9;data[879][7:5]<=3;data[879][4:0]<=3;
			data[880][11:8]<=6;data[880][7:5]<=3;data[880][4:0]<=2;
			data[881][11:8]<=9;data[881][7:5]<=3;data[881][4:0]<=16;
			data[882][11:8]<=0;data[882][7:5]<=4;data[882][4:0]<=4;
			data[883][11:8]<=9;data[883][7:5]<=3;data[883][4:0]<=2;
			data[884][11:8]<=11;data[884][7:5]<=3;data[884][4:0]<=2;
			data[885][11:8]<=9;data[885][7:5]<=3;data[885][4:0]<=3;
			data[886][11:8]<=6;data[886][7:5]<=3;data[886][4:0]<=2;
			data[887][11:8]<=9;data[887][7:5]<=3;data[887][4:0]<=3;
			data[888][11:8]<=2;data[888][7:5]<=3;data[888][4:0]<=4;
			data[889][11:8]<=2;data[889][7:5]<=3;data[889][4:0]<=2;
			data[890][11:8]<=4;data[890][7:5]<=3;data[890][4:0]<=2;
			data[891][11:8]<=6;data[891][7:5]<=3;data[891][4:0]<=2;
			data[892][11:8]<=11;data[892][7:5]<=3;data[892][4:0]<=2;
			data[893][11:8]<=2;data[893][7:5]<=3;data[893][4:0]<=4;
			data[894][11:8]<=6;data[894][7:5]<=3;data[894][4:0]<=2;
			data[895][11:8]<=9;data[895][7:5]<=3;data[895][4:0]<=2;
			data[896][11:8]<=4;data[896][7:5]<=2;data[896][4:0]<=8;
			data[897][11:8]<=9;data[897][7:5]<=3;data[897][4:0]<=8;
			data[898][11:8]<=0;data[898][7:5]<=4;data[898][4:0]<=4;
			data[899][11:8]<=0;data[899][7:5]<=4;data[899][4:0]<=4;
			data[900][11:8]<=9;data[900][7:5]<=4;data[900][4:0]<=4;
			data[901][11:8]<=11;data[901][7:5]<=4;data[901][4:0]<=4;
			data[902][11:8]<=2;data[902][7:5]<=3;data[902][4:0]<=4;
			data[903][11:8]<=4;data[903][7:5]<=3;data[903][4:0]<=2;
			data[904][11:8]<=9;data[904][7:5]<=4;data[904][4:0]<=2;
			data[905][11:8]<=9;data[905][7:5]<=4;data[905][4:0]<=4;
			data[906][11:8]<=11;data[906][7:5]<=4;data[906][4:0]<=4;
			data[907][11:8]<=2;data[907][7:5]<=3;data[907][4:0]<=2;
			data[908][11:8]<=4;data[908][7:5]<=3;data[908][4:0]<=2;
			data[909][11:8]<=9;data[909][7:5]<=4;data[909][4:0]<=4;
			data[910][11:8]<=6;data[910][7:5]<=3;data[910][4:0]<=4;
			data[911][11:8]<=4;data[911][7:5]<=3;data[911][4:0]<=4;
			data[912][11:8]<=4;data[912][7:5]<=3;data[912][4:0]<=4;
			data[913][11:8]<=2;data[913][7:5]<=3;data[913][4:0]<=2;
			data[914][11:8]<=13;data[914][7:5]<=4;data[914][4:0]<=2;
			data[915][11:8]<=13;data[915][7:5]<=4;data[915][4:0]<=4;
			data[916][11:8]<=2;data[916][7:5]<=3;data[916][4:0]<=4;
			data[917][11:8]<=13;data[917][7:5]<=4;data[917][4:0]<=4;
			data[918][11:8]<=9;data[918][7:5]<=4;data[918][4:0]<=4;
			data[919][11:8]<=9;data[919][7:5]<=4;data[919][4:0]<=4;
			data[920][11:8]<=11;data[920][7:5]<=4;data[920][4:0]<=4;
			data[921][11:8]<=2;data[921][7:5]<=3;data[921][4:0]<=4;
			data[922][11:8]<=4;data[922][7:5]<=3;data[922][4:0]<=2;
			data[923][11:8]<=9;data[923][7:5]<=4;data[923][4:0]<=2;
			data[924][11:8]<=9;data[924][7:5]<=4;data[924][4:0]<=4;
			data[925][11:8]<=11;data[925][7:5]<=4;data[925][4:0]<=4;
			data[926][11:8]<=2;data[926][7:5]<=3;data[926][4:0]<=2;
			data[927][11:8]<=4;data[927][7:5]<=3;data[927][4:0]<=2;
			data[928][11:8]<=9;data[928][7:5]<=4;data[928][4:0]<=4;
			data[929][11:8]<=6;data[929][7:5]<=3;data[929][4:0]<=4;
			data[930][11:8]<=4;data[930][7:5]<=3;data[930][4:0]<=4;
			data[931][11:8]<=2;data[931][7:5]<=3;data[931][4:0]<=2;
			data[932][11:8]<=13;data[932][7:5]<=4;data[932][4:0]<=2;
			data[933][11:8]<=13;data[933][7:5]<=4;data[933][4:0]<=4;
			data[934][11:8]<=2;data[934][7:5]<=3;data[934][4:0]<=12;

		end
		else if(wen_c)
			data[addr_c] <= data_c;
	end
	assign q_a = data[addr_a];
	assign q_b = data[addr_b];
	endmodule
